	component unsaved is
	end component unsaved;

	u0 : component unsaved
		port map (
		);

